`timescale 1ns/1ps

// Dual-port twiddle ROM for N=256 Kyber-style NTT over q=3329.
// Stores omega^i in Montgomery domain (value * R mod q, R=2^16 mod q).
module ntt_twiddle_rom # (
    parameter int WIDTH = 16,
    parameter int DEPTH = 256,
    parameter int ADDR_W = $clog2(DEPTH)
) (
    input  logic                 clk,
    input  logic                 en_a,
    input  logic [ADDR_W-1:0]    addr_a,
    output logic [WIDTH-1:0]     dout_a,
    input  logic                 en_b,
    input  logic [ADDR_W-1:0]    addr_b,
    output logic [WIDTH-1:0]     dout_b
);
    logic [WIDTH-1:0] rom [0:DEPTH-1];

    initial begin
        rom[0] = 16'd2285;
        rom[1] = 16'd2226;
        rom[2] = 16'd1223;
        rom[3] = 16'd817;
        rom[4] = 16'd573;
        rom[5] = 16'd3083;
        rom[6] = 16'd2476;
        rom[7] = 16'd2144;
        rom[8] = 16'd3158;
        rom[9] = 16'd422;
        rom[10] = 16'd516;
        rom[11] = 16'd2114;
        rom[12] = 16'd2648;
        rom[13] = 16'd1739;
        rom[14] = 16'd2931;
        rom[15] = 16'd3221;
        rom[16] = 16'd1493;
        rom[17] = 16'd2078;
        rom[18] = 16'd2036;
        rom[19] = 16'd1322;
        rom[20] = 16'd2500;
        rom[21] = 16'd2552;
        rom[22] = 16'd107;
        rom[23] = 16'd1819;
        rom[24] = 16'd962;
        rom[25] = 16'd3038;
        rom[26] = 16'd1711;
        rom[27] = 16'd2455;
        rom[28] = 16'd1787;
        rom[29] = 16'd418;
        rom[30] = 16'd448;
        rom[31] = 16'd958;
        rom[32] = 16'd2970;
        rom[33] = 16'd555;
        rom[34] = 16'd2777;
        rom[35] = 16'd603;
        rom[36] = 16'd264;
        rom[37] = 16'd1159;
        rom[38] = 16'd3058;
        rom[39] = 16'd2051;
        rom[40] = 16'd1577;
        rom[41] = 16'd177;
        rom[42] = 16'd3009;
        rom[43] = 16'd1218;
        rom[44] = 16'd732;
        rom[45] = 16'd2457;
        rom[46] = 16'd1821;
        rom[47] = 16'd996;
        rom[48] = 16'd287;
        rom[49] = 16'd1550;
        rom[50] = 16'd3047;
        rom[51] = 16'd1864;
        rom[52] = 16'd1727;
        rom[53] = 16'd2727;
        rom[54] = 16'd3082;
        rom[55] = 16'd2459;
        rom[56] = 16'd1855;
        rom[57] = 16'd1574;
        rom[58] = 16'd126;
        rom[59] = 16'd2142;
        rom[60] = 16'd3124;
        rom[61] = 16'd3173;
        rom[62] = 16'd677;
        rom[63] = 16'd1522;
        rom[64] = 16'd2571;
        rom[65] = 16'd430;
        rom[66] = 16'd652;
        rom[67] = 16'd1097;
        rom[68] = 16'd2004;
        rom[69] = 16'd778;
        rom[70] = 16'd3239;
        rom[71] = 16'd1799;
        rom[72] = 16'd622;
        rom[73] = 16'd587;
        rom[74] = 16'd3321;
        rom[75] = 16'd3193;
        rom[76] = 16'd1017;
        rom[77] = 16'd644;
        rom[78] = 16'd961;
        rom[79] = 16'd3021;
        rom[80] = 16'd1422;
        rom[81] = 16'd871;
        rom[82] = 16'd1491;
        rom[83] = 16'd2044;
        rom[84] = 16'd1458;
        rom[85] = 16'd1483;
        rom[86] = 16'd1908;
        rom[87] = 16'd2475;
        rom[88] = 16'd2127;
        rom[89] = 16'd2869;
        rom[90] = 16'd2167;
        rom[91] = 16'd220;
        rom[92] = 16'd411;
        rom[93] = 16'd329;
        rom[94] = 16'd2264;
        rom[95] = 16'd1869;
        rom[96] = 16'd1812;
        rom[97] = 16'd843;
        rom[98] = 16'd1015;
        rom[99] = 16'd610;
        rom[100] = 16'd383;
        rom[101] = 16'd3182;
        rom[102] = 16'd830;
        rom[103] = 16'd794;
        rom[104] = 16'd182;
        rom[105] = 16'd3094;
        rom[106] = 16'd2663;
        rom[107] = 16'd1994;
        rom[108] = 16'd608;
        rom[109] = 16'd349;
        rom[110] = 16'd2604;
        rom[111] = 16'd991;
        rom[112] = 16'd202;
        rom[113] = 16'd105;
        rom[114] = 16'd1785;
        rom[115] = 16'd384;
        rom[116] = 16'd3199;
        rom[117] = 16'd1119;
        rom[118] = 16'd2378;
        rom[119] = 16'd478;
        rom[120] = 16'd1468;
        rom[121] = 16'd1653;
        rom[122] = 16'd1469;
        rom[123] = 16'd1670;
        rom[124] = 16'd1758;
        rom[125] = 16'd3254;
        rom[126] = 16'd2054;
        rom[127] = 16'd1628;
        rom[128] = 16'd1044;
        rom[129] = 16'd1103;
        rom[130] = 16'd2106;
        rom[131] = 16'd2512;
        rom[132] = 16'd2756;
        rom[133] = 16'd246;
        rom[134] = 16'd853;
        rom[135] = 16'd1185;
        rom[136] = 16'd171;
        rom[137] = 16'd2907;
        rom[138] = 16'd2813;
        rom[139] = 16'd1215;
        rom[140] = 16'd681;
        rom[141] = 16'd1590;
        rom[142] = 16'd398;
        rom[143] = 16'd108;
        rom[144] = 16'd1836;
        rom[145] = 16'd1251;
        rom[146] = 16'd1293;
        rom[147] = 16'd2007;
        rom[148] = 16'd829;
        rom[149] = 16'd777;
        rom[150] = 16'd3222;
        rom[151] = 16'd1510;
        rom[152] = 16'd2367;
        rom[153] = 16'd291;
        rom[154] = 16'd1618;
        rom[155] = 16'd874;
        rom[156] = 16'd1542;
        rom[157] = 16'd2911;
        rom[158] = 16'd2881;
        rom[159] = 16'd2371;
        rom[160] = 16'd359;
        rom[161] = 16'd2774;
        rom[162] = 16'd552;
        rom[163] = 16'd2726;
        rom[164] = 16'd3065;
        rom[165] = 16'd2170;
        rom[166] = 16'd271;
        rom[167] = 16'd1278;
        rom[168] = 16'd1752;
        rom[169] = 16'd3152;
        rom[170] = 16'd320;
        rom[171] = 16'd2111;
        rom[172] = 16'd2597;
        rom[173] = 16'd872;
        rom[174] = 16'd1508;
        rom[175] = 16'd2333;
        rom[176] = 16'd3042;
        rom[177] = 16'd1779;
        rom[178] = 16'd282;
        rom[179] = 16'd1465;
        rom[180] = 16'd1602;
        rom[181] = 16'd602;
        rom[182] = 16'd247;
        rom[183] = 16'd870;
        rom[184] = 16'd1474;
        rom[185] = 16'd1755;
        rom[186] = 16'd3203;
        rom[187] = 16'd1187;
        rom[188] = 16'd205;
        rom[189] = 16'd156;
        rom[190] = 16'd2652;
        rom[191] = 16'd1807;
        rom[192] = 16'd758;
        rom[193] = 16'd2899;
        rom[194] = 16'd2677;
        rom[195] = 16'd2232;
        rom[196] = 16'd1325;
        rom[197] = 16'd2551;
        rom[198] = 16'd90;
        rom[199] = 16'd1530;
        rom[200] = 16'd2707;
        rom[201] = 16'd2742;
        rom[202] = 16'd8;
        rom[203] = 16'd136;
        rom[204] = 16'd2312;
        rom[205] = 16'd2685;
        rom[206] = 16'd2368;
        rom[207] = 16'd308;
        rom[208] = 16'd1907;
        rom[209] = 16'd2458;
        rom[210] = 16'd1838;
        rom[211] = 16'd1285;
        rom[212] = 16'd1871;
        rom[213] = 16'd1846;
        rom[214] = 16'd1421;
        rom[215] = 16'd854;
        rom[216] = 16'd1202;
        rom[217] = 16'd460;
        rom[218] = 16'd1162;
        rom[219] = 16'd3109;
        rom[220] = 16'd2918;
        rom[221] = 16'd3000;
        rom[222] = 16'd1065;
        rom[223] = 16'd1460;
        rom[224] = 16'd1517;
        rom[225] = 16'd2486;
        rom[226] = 16'd2314;
        rom[227] = 16'd2719;
        rom[228] = 16'd2946;
        rom[229] = 16'd147;
        rom[230] = 16'd2499;
        rom[231] = 16'd2535;
        rom[232] = 16'd3147;
        rom[233] = 16'd235;
        rom[234] = 16'd666;
        rom[235] = 16'd1335;
        rom[236] = 16'd2721;
        rom[237] = 16'd2980;
        rom[238] = 16'd725;
        rom[239] = 16'd2338;
        rom[240] = 16'd3127;
        rom[241] = 16'd3224;
        rom[242] = 16'd1544;
        rom[243] = 16'd2945;
        rom[244] = 16'd130;
        rom[245] = 16'd2210;
        rom[246] = 16'd951;
        rom[247] = 16'd2851;
        rom[248] = 16'd1861;
        rom[249] = 16'd1676;
        rom[250] = 16'd1860;
        rom[251] = 16'd1659;
        rom[252] = 16'd1571;
        rom[253] = 16'd75;
        rom[254] = 16'd1275;
        rom[255] = 16'd1701;
    end

    always_ff @(posedge clk) begin
        if (en_a) begin
            dout_a <= rom[addr_a];
        end
        if (en_b) begin
            dout_b <= rom[addr_b];
        end
    end

    // ROM-address safety assertions for an 8-stage (log2(256)) NTT fold.
    property p_addr_a_in_range;
        @(posedge clk) en_a |-> (addr_a < DEPTH);
    endproperty
    property p_addr_b_in_range;
        @(posedge clk) en_b |-> (addr_b < DEPTH);
    endproperty
    assert property (p_addr_a_in_range) else $fatal(1, "Twiddle ROM port A out-of-range access");
    assert property (p_addr_b_in_range) else $fatal(1, "Twiddle ROM port B out-of-range access");
endmodule
